module tlc_tb
